library verilog;
use verilog.vl_types.all;
entity output_encoder_vlg_vec_tst is
end output_encoder_vlg_vec_tst;
